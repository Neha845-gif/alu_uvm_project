`define width 8
`define no_of_transactions 5000
