package my_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "defines.sv"
    `include "seq_item.sv"
    `include "my_sequence.sv"
    `include "my_sequencer.sv"
    `include "my_driver.sv"
    `include "my_monitor.sv"
    `include "my_agent.sv"
    `include "my_scoreboard.sv"
    `include "my_coverage.sv"
    `include "my_env.sv"
    `include "my_test.sv"
endpackage
